
`ifndef ___uvm_apb_test__svh___
`define ___uvm_apb_test__svh___


   `include "test/uvm_apb_scoreboard.svh"           
   `include "test/uvm_apb_env.svh"                
   `include "test/uvm_apb_test.svh"               

// `include "uvm_apb_virtual_sequencer.svh"  
// `include "uvm_apb_virtual_sequence.svh"   

`endif
