`ifndef ___UVM_RESET_AGENT_SVH__
`define ___UVM_RESET_AGENT_SVH__


   `include "include/agent/reset_interface.svh"


   `include "include/agent/uvm_reset_sequence_item.svh"       
                                              
   `include "include/agent/uvm_reset_monitor.svh"             
                                              
   `include "include/agent/uvm_reset_driver.svh"       
   `include "include/agent/uvm_reset_sequencer.svh"    
   `include "include/agent/uvm_reset_agent.svh"        

   `include "include/sequence/uvm_reset_sequence.svh"    
                                              
`endif
