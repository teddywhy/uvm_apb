`ifndef ___uvm_reset_agent__svh___
`define ___uvm_reset_agent__svh___


   `include "agent/reset_interface.svh"


   `include "agent/uvm_reset_sequence_item.svh"       
                                      
   `include "agent/uvm_reset_monitor.svh"             
                                      
   `include "agent/uvm_reset_driver.svh"       
   `include "agent/uvm_reset_sequencer.svh"    
   `include "agent/uvm_reset_agent.svh"        

   `include "sequence/uvm_reset_sequence.svh"    
                                              
`endif
