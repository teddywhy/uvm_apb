`ifndef ____uvm_apb__svh____
`define ____uvm_apb__svh____

   `include "agent/apb_parameter.svh"
   `include "agent/apb_interface.svh"


   `include "agent/uvm_apb_sequence_item.svh"       
                              
   `include "agent/uvm_apb_monitor.svh"             
   `include "agent/uvm_apb_request_monitor.svh"             
                              
   `include "agent/uvm_apb_master_driver.svh"       
   `include "agent/uvm_apb_master_sequencer.svh"    
   `include "agent/uvm_apb_master_agent.svh"        
                              
   `include "agent/uvm_apb_slave_driver.svh"        
   `include "agent/uvm_apb_slave_sequencer.svh"     
   `include "agent/uvm_apb_slave_agent.svh"         

   `include "sequence/uvm_apb_slave_response_sequence.svh"

   `include "sequence/uvm_apb_master_sequence.svh"
   `include "sequence/uvm_apb_master_sequence_r.svh"
   `include "sequence/uvm_apb_master_sequence_w.svh"

`endif


