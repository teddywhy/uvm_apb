
`ifndef ___UVM_APB_TEST_SVH__
`define ___UVM_APB_TEST_SVH__

   `include "uvm_apb_test/uvm_apb_scoreboard.svh"           
   `include "uvm_apb_test/uvm_apb_env.svh"                
   `include "uvm_apb_test/uvm_apb_test.svh"               

// `include "uvm_apb_virtual_sequencer.svh"  
// `include "uvm_apb_virtual_sequence.svh"   

`endif
