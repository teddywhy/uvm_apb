`ifndef ___UVM_APB_AGENT_SVH__
`define ___UVM_APB_AGENT_SVH__

   `include "uvm_apb_agent/apb_parameter.svh"
   `include "uvm_apb_agent/apb_interface.svh"


   `include "uvm_apb_agent/uvm_apb_sequence_item.svh"       
                                              
   `include "uvm_apb_agent/uvm_apb_monitor.svh"             
   `include "uvm_apb_agent/uvm_apb_request_monitor.svh"             
                                              
   `include "uvm_apb_agent/uvm_apb_master_driver.svh"       
   `include "uvm_apb_agent/uvm_apb_master_sequencer.svh"    
   `include "uvm_apb_agent/uvm_apb_master_agent.svh"        
                                              
   `include "uvm_apb_agent/uvm_apb_slave_driver.svh"        
   `include "uvm_apb_agent/uvm_apb_slave_sequencer.svh"     
   `include "uvm_apb_agent/uvm_apb_slave_agent.svh"         

   `include "uvm_apb_agent/uvm_apb_slave_response_sequence.svh"

   `include "uvm_apb_agent/sequence/uvm_apb_master_sequence.svh"
   `include "uvm_apb_agent/sequence/uvm_apb_master_sequence_r.svh"
   `include "uvm_apb_agent/sequence/uvm_apb_master_sequence_w.svh"

`endif
