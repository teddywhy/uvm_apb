
package uvm_apb_master_test_pkg;
    
    import uvm_apb_agent_pkg::*;
    
    `include "uvm_apb_master_env.svh"
    `include "uvm_apb_master_scoreboard.svh"

    `include "uvm_apb_master_test.svh"

endpackage: uvm_apb_master_test_pkg     
