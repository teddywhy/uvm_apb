
`ifndef ___uvm_apb_master_test__svh___
`define ___uvm_apb_master_test__svh___

   `include "master_test/uvm_apb_master_scoreboard.svh"     
   `include "master_test/uvm_apb_master_env.svh"            
   `include "master_test/uvm_apb_master_test.svh"              

`endif
   