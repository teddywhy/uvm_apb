
 typedef struct packed
 {
   int unsigned   ADDR_WIDTH ;
   int unsigned   DATA_WIDTH ;
 }
 apb_parameter_t;

 parameter apb_parameter_t apb_parameter =
 '{
       ADDR_WIDTH : 11  ,
       DATA_WIDTH : 32
  };


