
`ifndef ___UVM_APB_MASTER_TEST_SVH__
`define ___UVM_APB_MASTER_TEST_SVH__

   `include "uvm_apb_master_test/uvm_apb_master_scoreboard.svh"
     
   `include "uvm_apb_master_test/uvm_apb_master_env.svh"
   `include "uvm_apb_master_test/uvm_apb_master_test.svh"
   
`endif
   