`ifndef ___UVM_RESET_AGENT_SVH__
`define ___UVM_RESET_AGENT_SVH__


   `include "uvm_reset_agent/reset_interface.svh"


   `include "uvm_reset_agent/uvm_reset_sequence_item.svh"       
                                              
   `include "uvm_reset_agent/uvm_reset_monitor.svh"             
                                              
   `include "uvm_reset_agent/uvm_reset_driver.svh"       
   `include "uvm_reset_agent/uvm_reset_sequencer.svh"    
   `include "uvm_reset_agent/uvm_reset_agent.svh"        

   `include "uvm_reset_agent/uvm_reset_sequence.svh"    
                                              
`endif
