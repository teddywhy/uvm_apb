
`ifndef ___UVM_APB_SEQUENCE_SVH__
`define ___UVM_APB_SEQUENCE_SVH__

   `include "uvm_apb_sequence/uvm_apb_master_sequence.svh"
   `include "uvm_apb_sequence/uvm_apb_master_sequence_r.svh"
   `include "uvm_apb_sequence/uvm_apb_master_sequence_w.svh"

`endif
