
 typedef struct packed
 {
   int unsigned   WIDTH ;
 }
 reset_parameter_t;

 parameter reset_parameter_t reset_parameter =
 '{
       WIDTH : 8 
  };


