
package uvm_apb_sequence_pkg;

  `include "uvm_apb_sequence.svh"
  `include "uvm_apb_sequence_r.svh"
  `include "uvm_apb_sequence_w.svh"

endpackage : uvm_apb_sequence_pkg