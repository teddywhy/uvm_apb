


package uvm_apb_package;


// `include "include/agent/apb_parameter.svh"
// `include "include/agent/apb_interface.svh"


   `include "include/agent/uvm_apb_sequence_item.svh"       
                                      
   `include "include/agent/uvm_apb_monitor.svh"             
   `include "include/agent/uvm_apb_request_monitor.svh"             
                                      
   `include "include/agent/uvm_apb_master_driver.svh"       
   `include "include/agent/uvm_apb_master_sequencer.svh"    
   `include "include/agent/uvm_apb_master_agent.svh"        
                                      
   `include "include/agent/uvm_apb_slave_driver.svh"        
   `include "include/agent/uvm_apb_slave_sequencer.svh"     
   `include "include/agent/uvm_apb_slave_agent.svh"         

   `include "include/sequence/uvm_apb_slave_response_sequence.svh"

   `include "include/sequence/uvm_apb_master_sequence.svh"
   `include "include/sequence/uvm_apb_master_sequence_r.svh"
   `include "include/sequence/uvm_apb_master_sequence_w.svh"

endpackage: uvm_apb_package     
